/*
 Produced by NSL Core(version=20140126), IP ARCH, Inc. Sun Aug 14 20:41:10 2016
 Licensed to :EVALUATION USER
*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module duty2 ( p_reset , m_clock , Vin , dnum , V0 , setduty , exec );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input [3:0] Vin;
  wire [3:0] Vin;
  input [1:0] dnum;
  wire [1:0] dnum;
  output [3:0] V0;
  wire [3:0] V0;
  input setduty;
  wire setduty;
  input exec;
  wire exec;
  reg [5:0] cnt;
  reg [1:0] d;
  wire _net_0;
  wire _net_1;
  wire _net_2;
  wire _net_3;
  wire _net_4;
  wire _net_5;
  wire _net_6;
  wire _net_7;
  wire _net_8;
  wire _net_9;
  wire _net_10;
  wire _net_11;
  wire _net_12;
  wire _net_13;
  wire _net_14;
  wire _net_15;
  wire _net_16;
  wire _net_17;
  wire _net_18;
  wire _net_19;
  wire _net_20;
  wire _net_21;
  wire _net_22;
  wire _net_23;
  wire _net_24;
  wire _net_25;
  wire _net_26;
  wire _net_27;
  wire _net_28;
  wire _net_29;
  wire _net_30;
  wire _net_31;
  wire _net_32;
  wire _net_33;
  wire _net_34;
  wire _net_35;
  wire _net_36;
  wire _net_37;
  wire _net_38;
  wire _net_39;
  wire _net_40;
  wire _net_41;
  wire _net_42;
  wire _net_43;
  wire _net_44;
  wire _net_45;
  wire _net_46;
  wire _net_47;
  wire _net_48;
  wire _net_49;
  wire _net_50;
  wire _net_51;
  wire _net_52;
  wire _net_53;
  wire _net_54;
  wire _net_55;
  wire _net_56;
  wire _net_57;
  wire _net_58;
  wire _net_59;
  wire _net_60;
  wire _net_61;
  wire _net_62;
  wire _net_63;
  wire _net_64;
  wire _net_65;
  wire _net_66;
  wire _net_67;
  wire _net_68;
  wire _net_69;
  wire _net_70;
  wire _net_71;
  wire _net_72;
  wire _net_73;
  wire _net_74;
  wire _net_75;
  wire _net_76;
  wire _net_77;
  wire _net_78;
  wire _net_79;
  wire _net_80;
  wire _net_81;
  wire _net_82;
  wire _net_83;
  wire _net_84;
  wire _net_85;
  wire _net_86;
  wire _net_87;
  wire _net_88;
  wire _net_89;
  wire _net_90;
  wire _net_91;
  wire _net_92;
  wire _net_93;
  wire _net_94;
  wire _net_95;
  wire _net_96;
  wire _net_97;
  wire _net_98;
  wire _net_99;
  wire _net_100;
  wire _net_101;
  wire _net_102;
  wire _net_103;
  wire _net_104;
  wire _net_105;
  wire _net_106;
  wire _net_107;
  wire _net_108;
  wire _net_109;
  wire _net_110;
  wire _net_111;
  wire _net_112;
  wire _net_113;
  wire _net_114;
  wire _net_115;
  wire _net_116;
  wire _net_117;
  wire _net_118;
  wire _net_119;
  wire _net_120;
  wire _net_121;
  wire _net_122;
  wire _net_123;
  wire _net_124;
  wire _net_125;
  wire _net_126;
  wire _net_127;
  wire _net_128;
  wire _net_129;
  wire _net_130;
  wire _net_131;
  wire _net_132;
  wire _net_133;

   assign  _net_0 = 
// synthesis translate_off
// synopsys translate_off
(exec)? 
// synthesis translate_on
// synopsys translate_on
((exec)?(cnt != 6'b011111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_1 = 
// synthesis translate_off
// synopsys translate_off
(exec)? 
// synthesis translate_on
// synopsys translate_on
((exec)?(cnt==6'b011111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_2 = (d==2'b00);
   assign  _net_3 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_4 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_5 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_6 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_7 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_8 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_9 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_10 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b011000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_11 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_12 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_13 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_14 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_15 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_16 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_17 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_18 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b010000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_19 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_20 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_21 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_22 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_23 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_24 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_25 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_26 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b001000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_27 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_28 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_29 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_30 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_31 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_32 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_33 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_34 = 
// synthesis translate_off
// synopsys translate_off
(_net_2)? 
// synthesis translate_on
// synopsys translate_on
((_net_2)?(cnt==6'b000000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_35 = (d==2'b01);
   assign  _net_36 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_37 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_38 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_39 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_40 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_41 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_42 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_43 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b011000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_44 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_45 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_46 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_47 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_48 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_49 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_50 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_51 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b010000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_52 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_53 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_54 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_55 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_56 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_57 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_58 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_59 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b001000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_60 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_61 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_62 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_63 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_64 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_65 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_66 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_67 = 
// synthesis translate_off
// synopsys translate_off
(_net_35)? 
// synthesis translate_on
// synopsys translate_on
((_net_35)?(cnt==6'b000000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_68 = (d==2'b10);
   assign  _net_69 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_70 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_71 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_72 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_73 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_74 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_75 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_76 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b011000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_77 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_78 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_79 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_80 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_81 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_82 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_83 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_84 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b010000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_85 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_86 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_87 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_88 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_89 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_90 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_91 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_92 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b001000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_93 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_94 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_95 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_96 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_97 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_98 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_99 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_100 = 
// synthesis translate_off
// synopsys translate_off
(_net_68)? 
// synthesis translate_on
// synopsys translate_on
((_net_68)?(cnt==6'b000000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_101 = (d==2'b11);
   assign  _net_102 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_103 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_104 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_105 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_106 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_107 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_108 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_109 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b011000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_110 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_111 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_112 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_113 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_114 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_115 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_116 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_117 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b010000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_118 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_119 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_120 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_121 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_122 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_123 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_124 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_125 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b001000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_126 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000111):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_127 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000110):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_128 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000101):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_129 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000100):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_130 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000011):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_131 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000010):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_132 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000001):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_133 = 
// synthesis translate_off
// synopsys translate_off
(_net_101)? 
// synthesis translate_on
// synopsys translate_on
((_net_101)?(cnt==6'b000000):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)&(_net_101&_net_132))|(((_net_101&_net_133)|(_net_101&_net_132))&(_net_101&_net_131)))|((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))&(_net_101&_net_130)))|(((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))&(_net_101&_net_129)))|((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))&(_net_101&_net_128)))|(((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))&(_net_101&_net_127)))|((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))&(_net_101&_net_126)))|(((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))&(_net_101&_net_125)))|((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))&(_net_101&_net_124)))|(((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))&(_net_101&_net_123)))|((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))&(_net_101&_net_122)))|(((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))&(_net_101&_net_121)))|((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))&(_net_101&_net_120)))|(((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))&(_net_101&_net_119)))|((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))&(_net_101&_net_118)))|(((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))&(_net_101&_net_117)))|((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))&(_net_101&_net_116)))|(((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))&(_net_101&_net_115)))|((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))&(_net_101&_net_114)))|(((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))&(_net_101&_net_113)))|((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))&(_net_101&_net_112)))|(((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))&(_net_101&_net_111)))|((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))&(_net_101&_net_110)))|(((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))&(_net_101&_net_109)))|((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))&(_net_101&_net_108)))|(((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))&(_net_101&_net_107)))|((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))&(_net_101&_net_106)))|(((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))&(_net_101&_net_105)))|((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))&(_net_101&_net_104)))|(((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))&(_net_101&_net_103)))|((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))&(_net_101&_net_102)))|(((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))&(_net_68&_net_100)))|((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))&(_net_68&_net_99)))|(((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))&(_net_68&_net_98)))|((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))&(_net_68&_net_97)))|(((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))&(_net_68&_net_96)))|((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))&(_net_68&_net_95)))|(((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))&(_net_68&_net_94)))|((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))&(_net_68&_net_93)))|(((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))&(_net_68&_net_92)))|((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))&(_net_68&_net_91)))|(((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))&(_net_68&_net_90)))|((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))&(_net_68&_net_89)))|(((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))&(_net_68&_net_88)))|((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))&(_net_68&_net_87)))|(((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))&(_net_68&_net_86)))|((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))&(_net_68&_net_85)))|(((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))&(_net_68&_net_84)))|((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))&(_net_68&_net_83)))|(((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))&(_net_68&_net_82)))|((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))&(_net_68&_net_81)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))&(_net_68&_net_80)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))&(_net_68&_net_79)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))&(_net_68&_net_78)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))&(_net_68&_net_77)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))&(_net_68&_net_76)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))&(_net_68&_net_75)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))&(_net_68&_net_74)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))&(_net_68&_net_73)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))&(_net_68&_net_72)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))&(_net_68&_net_71)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))&(_net_68&_net_70)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))&(_net_68&_net_69)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))&(_net_35&_net_67)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))&(_net_35&_net_66)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))&(_net_35&_net_65)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))&(_net_35&_net_64)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))&(_net_35&_net_63)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))&(_net_35&_net_62)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))&(_net_35&_net_61)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))&(_net_35&_net_60)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))&(_net_35&_net_59)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))&(_net_35&_net_58)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))&(_net_35&_net_57)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))&(_net_35&_net_56)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))&(_net_35&_net_55)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))&(_net_35&_net_54)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))&(_net_35&_net_53)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))&(_net_35&_net_52)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))&(_net_35&_net_51)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))&(_net_35&_net_50)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))&(_net_35&_net_49)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))&(_net_35&_net_48)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))&(_net_35&_net_47)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))&(_net_35&_net_46)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))&(_net_35&_net_45)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))&(_net_35&_net_44)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))&(_net_35&_net_43)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))&(_net_35&_net_42)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))&(_net_35&_net_41)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))&(_net_35&_net_40)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))&(_net_35&_net_39)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))&(_net_35&_net_38)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))&(_net_35&_net_37)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))&(_net_35&_net_36)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))&(_net_2&_net_34)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))&(_net_2&_net_33)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))&(_net_2&_net_32)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))&(_net_2&_net_31)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))&(_net_2&_net_30)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))&(_net_2&_net_29)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))&(_net_2&_net_28)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))&(_net_2&_net_27)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))&(_net_2&_net_26)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))&(_net_2&_net_25)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))&(_net_2&_net_24)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))&(_net_2&_net_23)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))&(_net_2&_net_22)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))&(_net_2&_net_21)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))&(_net_2&_net_20)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))&(_net_2&_net_19)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))&(_net_2&_net_18)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))&(_net_2&_net_17)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))&(_net_2&_net_16)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))&(_net_2&_net_15)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))&(_net_2&_net_14)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))&(_net_2&_net_13)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))&(_net_2&_net_12)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))&(_net_2&_net_11)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))&(_net_2&_net_10)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))&(_net_2&_net_9)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))&(_net_2&_net_8)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))&(_net_2&_net_7)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))&(_net_2&_net_6)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))|(_net_2&_net_6))&(_net_2&_net_5)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))|(_net_2&_net_6))|(_net_2&_net_5))&(_net_2&_net_4)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))|(_net_2&_net_6))|(_net_2&_net_5))|(_net_2&_net_4))&(_net_2&_net_3))))
 begin $display("Warning: assign collision(duty2:V0) at %d",$time);
if ((_net_101&_net_133)) $display("assert ((_net_101&_net_133)) line 135 at %d\n",$time);
if ((_net_101&_net_132)) $display("assert ((_net_101&_net_132)) line 136 at %d\n",$time);
if ((_net_101&_net_131)) $display("assert ((_net_101&_net_131)) line 137 at %d\n",$time);
if ((_net_101&_net_130)) $display("assert ((_net_101&_net_130)) line 138 at %d\n",$time);
if ((_net_101&_net_129)) $display("assert ((_net_101&_net_129)) line 139 at %d\n",$time);
if ((_net_101&_net_128)) $display("assert ((_net_101&_net_128)) line 140 at %d\n",$time);
if ((_net_101&_net_127)) $display("assert ((_net_101&_net_127)) line 141 at %d\n",$time);
if ((_net_101&_net_126)) $display("assert ((_net_101&_net_126)) line 142 at %d\n",$time);
if ((_net_101&_net_125)) $display("assert ((_net_101&_net_125)) line 143 at %d\n",$time);
if ((_net_101&_net_124)) $display("assert ((_net_101&_net_124)) line 144 at %d\n",$time);
if ((_net_101&_net_123)) $display("assert ((_net_101&_net_123)) line 145 at %d\n",$time);
if ((_net_101&_net_122)) $display("assert ((_net_101&_net_122)) line 146 at %d\n",$time);
if ((_net_101&_net_121)) $display("assert ((_net_101&_net_121)) line 147 at %d\n",$time);
if ((_net_101&_net_120)) $display("assert ((_net_101&_net_120)) line 148 at %d\n",$time);
if ((_net_101&_net_119)) $display("assert ((_net_101&_net_119)) line 149 at %d\n",$time);
if ((_net_101&_net_118)) $display("assert ((_net_101&_net_118)) line 150 at %d\n",$time);
if ((_net_101&_net_117)) $display("assert ((_net_101&_net_117)) line 151 at %d\n",$time);
if ((_net_101&_net_116)) $display("assert ((_net_101&_net_116)) line 152 at %d\n",$time);
if ((_net_101&_net_115)) $display("assert ((_net_101&_net_115)) line 153 at %d\n",$time);
if ((_net_101&_net_114)) $display("assert ((_net_101&_net_114)) line 154 at %d\n",$time);
if ((_net_101&_net_113)) $display("assert ((_net_101&_net_113)) line 155 at %d\n",$time);
if ((_net_101&_net_112)) $display("assert ((_net_101&_net_112)) line 156 at %d\n",$time);
if ((_net_101&_net_111)) $display("assert ((_net_101&_net_111)) line 157 at %d\n",$time);
if ((_net_101&_net_110)) $display("assert ((_net_101&_net_110)) line 158 at %d\n",$time);
if ((_net_101&_net_109)) $display("assert ((_net_101&_net_109)) line 159 at %d\n",$time);
if ((_net_101&_net_108)) $display("assert ((_net_101&_net_108)) line 160 at %d\n",$time);
if ((_net_101&_net_107)) $display("assert ((_net_101&_net_107)) line 161 at %d\n",$time);
if ((_net_101&_net_106)) $display("assert ((_net_101&_net_106)) line 162 at %d\n",$time);
if ((_net_101&_net_105)) $display("assert ((_net_101&_net_105)) line 163 at %d\n",$time);
if ((_net_101&_net_104)) $display("assert ((_net_101&_net_104)) line 164 at %d\n",$time);
if ((_net_101&_net_103)) $display("assert ((_net_101&_net_103)) line 165 at %d\n",$time);
if ((_net_101&_net_102)) $display("assert ((_net_101&_net_102)) line 166 at %d\n",$time);
if ((_net_68&_net_100)) $display("assert ((_net_68&_net_100)) line 98 at %d\n",$time);
if ((_net_68&_net_99)) $display("assert ((_net_68&_net_99)) line 99 at %d\n",$time);
if ((_net_68&_net_98)) $display("assert ((_net_68&_net_98)) line 100 at %d\n",$time);
if ((_net_68&_net_97)) $display("assert ((_net_68&_net_97)) line 101 at %d\n",$time);
if ((_net_68&_net_96)) $display("assert ((_net_68&_net_96)) line 102 at %d\n",$time);
if ((_net_68&_net_95)) $display("assert ((_net_68&_net_95)) line 103 at %d\n",$time);
if ((_net_68&_net_94)) $display("assert ((_net_68&_net_94)) line 104 at %d\n",$time);
if ((_net_68&_net_93)) $display("assert ((_net_68&_net_93)) line 105 at %d\n",$time);
if ((_net_68&_net_92)) $display("assert ((_net_68&_net_92)) line 106 at %d\n",$time);
if ((_net_68&_net_91)) $display("assert ((_net_68&_net_91)) line 107 at %d\n",$time);
if ((_net_68&_net_90)) $display("assert ((_net_68&_net_90)) line 108 at %d\n",$time);
if ((_net_68&_net_89)) $display("assert ((_net_68&_net_89)) line 109 at %d\n",$time);
if ((_net_68&_net_88)) $display("assert ((_net_68&_net_88)) line 110 at %d\n",$time);
if ((_net_68&_net_87)) $display("assert ((_net_68&_net_87)) line 111 at %d\n",$time);
if ((_net_68&_net_86)) $display("assert ((_net_68&_net_86)) line 112 at %d\n",$time);
if ((_net_68&_net_85)) $display("assert ((_net_68&_net_85)) line 113 at %d\n",$time);
if ((_net_68&_net_84)) $display("assert ((_net_68&_net_84)) line 114 at %d\n",$time);
if ((_net_68&_net_83)) $display("assert ((_net_68&_net_83)) line 115 at %d\n",$time);
if ((_net_68&_net_82)) $display("assert ((_net_68&_net_82)) line 116 at %d\n",$time);
if ((_net_68&_net_81)) $display("assert ((_net_68&_net_81)) line 117 at %d\n",$time);
if ((_net_68&_net_80)) $display("assert ((_net_68&_net_80)) line 118 at %d\n",$time);
if ((_net_68&_net_79)) $display("assert ((_net_68&_net_79)) line 119 at %d\n",$time);
if ((_net_68&_net_78)) $display("assert ((_net_68&_net_78)) line 120 at %d\n",$time);
if ((_net_68&_net_77)) $display("assert ((_net_68&_net_77)) line 121 at %d\n",$time);
if ((_net_68&_net_76)) $display("assert ((_net_68&_net_76)) line 122 at %d\n",$time);
if ((_net_68&_net_75)) $display("assert ((_net_68&_net_75)) line 123 at %d\n",$time);
if ((_net_68&_net_74)) $display("assert ((_net_68&_net_74)) line 124 at %d\n",$time);
if ((_net_68&_net_73)) $display("assert ((_net_68&_net_73)) line 125 at %d\n",$time);
if ((_net_68&_net_72)) $display("assert ((_net_68&_net_72)) line 126 at %d\n",$time);
if ((_net_68&_net_71)) $display("assert ((_net_68&_net_71)) line 127 at %d\n",$time);
if ((_net_68&_net_70)) $display("assert ((_net_68&_net_70)) line 128 at %d\n",$time);
if ((_net_68&_net_69)) $display("assert ((_net_68&_net_69)) line 129 at %d\n",$time);
if ((_net_35&_net_67)) $display("assert ((_net_35&_net_67)) line 62 at %d\n",$time);
if ((_net_35&_net_66)) $display("assert ((_net_35&_net_66)) line 63 at %d\n",$time);
if ((_net_35&_net_65)) $display("assert ((_net_35&_net_65)) line 64 at %d\n",$time);
if ((_net_35&_net_64)) $display("assert ((_net_35&_net_64)) line 65 at %d\n",$time);
if ((_net_35&_net_63)) $display("assert ((_net_35&_net_63)) line 66 at %d\n",$time);
if ((_net_35&_net_62)) $display("assert ((_net_35&_net_62)) line 67 at %d\n",$time);
if ((_net_35&_net_61)) $display("assert ((_net_35&_net_61)) line 68 at %d\n",$time);
if ((_net_35&_net_60)) $display("assert ((_net_35&_net_60)) line 69 at %d\n",$time);
if ((_net_35&_net_59)) $display("assert ((_net_35&_net_59)) line 70 at %d\n",$time);
if ((_net_35&_net_58)) $display("assert ((_net_35&_net_58)) line 71 at %d\n",$time);
if ((_net_35&_net_57)) $display("assert ((_net_35&_net_57)) line 72 at %d\n",$time);
if ((_net_35&_net_56)) $display("assert ((_net_35&_net_56)) line 73 at %d\n",$time);
if ((_net_35&_net_55)) $display("assert ((_net_35&_net_55)) line 74 at %d\n",$time);
if ((_net_35&_net_54)) $display("assert ((_net_35&_net_54)) line 75 at %d\n",$time);
if ((_net_35&_net_53)) $display("assert ((_net_35&_net_53)) line 76 at %d\n",$time);
if ((_net_35&_net_52)) $display("assert ((_net_35&_net_52)) line 77 at %d\n",$time);
if ((_net_35&_net_51)) $display("assert ((_net_35&_net_51)) line 78 at %d\n",$time);
if ((_net_35&_net_50)) $display("assert ((_net_35&_net_50)) line 79 at %d\n",$time);
if ((_net_35&_net_49)) $display("assert ((_net_35&_net_49)) line 80 at %d\n",$time);
if ((_net_35&_net_48)) $display("assert ((_net_35&_net_48)) line 81 at %d\n",$time);
if ((_net_35&_net_47)) $display("assert ((_net_35&_net_47)) line 82 at %d\n",$time);
if ((_net_35&_net_46)) $display("assert ((_net_35&_net_46)) line 83 at %d\n",$time);
if ((_net_35&_net_45)) $display("assert ((_net_35&_net_45)) line 84 at %d\n",$time);
if ((_net_35&_net_44)) $display("assert ((_net_35&_net_44)) line 85 at %d\n",$time);
if ((_net_35&_net_43)) $display("assert ((_net_35&_net_43)) line 86 at %d\n",$time);
if ((_net_35&_net_42)) $display("assert ((_net_35&_net_42)) line 87 at %d\n",$time);
if ((_net_35&_net_41)) $display("assert ((_net_35&_net_41)) line 88 at %d\n",$time);
if ((_net_35&_net_40)) $display("assert ((_net_35&_net_40)) line 89 at %d\n",$time);
if ((_net_35&_net_39)) $display("assert ((_net_35&_net_39)) line 90 at %d\n",$time);
if ((_net_35&_net_38)) $display("assert ((_net_35&_net_38)) line 91 at %d\n",$time);
if ((_net_35&_net_37)) $display("assert ((_net_35&_net_37)) line 92 at %d\n",$time);
if ((_net_35&_net_36)) $display("assert ((_net_35&_net_36)) line 93 at %d\n",$time);
if ((_net_2&_net_34)) $display("assert ((_net_2&_net_34)) line 26 at %d\n",$time);
if ((_net_2&_net_33)) $display("assert ((_net_2&_net_33)) line 27 at %d\n",$time);
if ((_net_2&_net_32)) $display("assert ((_net_2&_net_32)) line 28 at %d\n",$time);
if ((_net_2&_net_31)) $display("assert ((_net_2&_net_31)) line 29 at %d\n",$time);
if ((_net_2&_net_30)) $display("assert ((_net_2&_net_30)) line 30 at %d\n",$time);
if ((_net_2&_net_29)) $display("assert ((_net_2&_net_29)) line 31 at %d\n",$time);
if ((_net_2&_net_28)) $display("assert ((_net_2&_net_28)) line 32 at %d\n",$time);
if ((_net_2&_net_27)) $display("assert ((_net_2&_net_27)) line 33 at %d\n",$time);
if ((_net_2&_net_26)) $display("assert ((_net_2&_net_26)) line 34 at %d\n",$time);
if ((_net_2&_net_25)) $display("assert ((_net_2&_net_25)) line 35 at %d\n",$time);
if ((_net_2&_net_24)) $display("assert ((_net_2&_net_24)) line 36 at %d\n",$time);
if ((_net_2&_net_23)) $display("assert ((_net_2&_net_23)) line 37 at %d\n",$time);
if ((_net_2&_net_22)) $display("assert ((_net_2&_net_22)) line 38 at %d\n",$time);
if ((_net_2&_net_21)) $display("assert ((_net_2&_net_21)) line 39 at %d\n",$time);
if ((_net_2&_net_20)) $display("assert ((_net_2&_net_20)) line 40 at %d\n",$time);
if ((_net_2&_net_19)) $display("assert ((_net_2&_net_19)) line 41 at %d\n",$time);
if ((_net_2&_net_18)) $display("assert ((_net_2&_net_18)) line 42 at %d\n",$time);
if ((_net_2&_net_17)) $display("assert ((_net_2&_net_17)) line 43 at %d\n",$time);
if ((_net_2&_net_16)) $display("assert ((_net_2&_net_16)) line 44 at %d\n",$time);
if ((_net_2&_net_15)) $display("assert ((_net_2&_net_15)) line 45 at %d\n",$time);
if ((_net_2&_net_14)) $display("assert ((_net_2&_net_14)) line 46 at %d\n",$time);
if ((_net_2&_net_13)) $display("assert ((_net_2&_net_13)) line 47 at %d\n",$time);
if ((_net_2&_net_12)) $display("assert ((_net_2&_net_12)) line 48 at %d\n",$time);
if ((_net_2&_net_11)) $display("assert ((_net_2&_net_11)) line 49 at %d\n",$time);
if ((_net_2&_net_10)) $display("assert ((_net_2&_net_10)) line 50 at %d\n",$time);
if ((_net_2&_net_9)) $display("assert ((_net_2&_net_9)) line 51 at %d\n",$time);
if ((_net_2&_net_8)) $display("assert ((_net_2&_net_8)) line 52 at %d\n",$time);
if ((_net_2&_net_7)) $display("assert ((_net_2&_net_7)) line 53 at %d\n",$time);
if ((_net_2&_net_6)) $display("assert ((_net_2&_net_6)) line 54 at %d\n",$time);
if ((_net_2&_net_5)) $display("assert ((_net_2&_net_5)) line 55 at %d\n",$time);
if ((_net_2&_net_4)) $display("assert ((_net_2&_net_4)) line 56 at %d\n",$time);
if ((_net_2&_net_3)) $display("assert ((_net_2&_net_3)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  V0 = 
// synthesis translate_off
// synopsys translate_off
(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)&(_net_101&_net_132))|(((_net_101&_net_133)|(_net_101&_net_132))&(_net_101&_net_131)))|((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))&(_net_101&_net_130)))|(((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))&(_net_101&_net_129)))|((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))&(_net_101&_net_128)))|(((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))&(_net_101&_net_127)))|((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))&(_net_101&_net_126)))|(((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))&(_net_101&_net_125)))|((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))&(_net_101&_net_124)))|(((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))&(_net_101&_net_123)))|((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))&(_net_101&_net_122)))|(((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))&(_net_101&_net_121)))|((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))&(_net_101&_net_120)))|(((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))&(_net_101&_net_119)))|((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))&(_net_101&_net_118)))|(((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))&(_net_101&_net_117)))|((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))&(_net_101&_net_116)))|(((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))&(_net_101&_net_115)))|((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))&(_net_101&_net_114)))|(((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))&(_net_101&_net_113)))|((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))&(_net_101&_net_112)))|(((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))&(_net_101&_net_111)))|((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))&(_net_101&_net_110)))|(((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))&(_net_101&_net_109)))|((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))&(_net_101&_net_108)))|(((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))&(_net_101&_net_107)))|((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))&(_net_101&_net_106)))|(((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))&(_net_101&_net_105)))|((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))&(_net_101&_net_104)))|(((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))&(_net_101&_net_103)))|((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))&(_net_101&_net_102)))|(((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))&(_net_68&_net_100)))|((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))&(_net_68&_net_99)))|(((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))&(_net_68&_net_98)))|((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))&(_net_68&_net_97)))|(((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))&(_net_68&_net_96)))|((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))&(_net_68&_net_95)))|(((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))&(_net_68&_net_94)))|((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))&(_net_68&_net_93)))|(((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))&(_net_68&_net_92)))|((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))&(_net_68&_net_91)))|(((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))&(_net_68&_net_90)))|((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))&(_net_68&_net_89)))|(((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))&(_net_68&_net_88)))|((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))&(_net_68&_net_87)))|(((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))&(_net_68&_net_86)))|((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))&(_net_68&_net_85)))|(((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))&(_net_68&_net_84)))|((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))&(_net_68&_net_83)))|(((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))&(_net_68&_net_82)))|((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))&(_net_68&_net_81)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))&(_net_68&_net_80)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))&(_net_68&_net_79)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))&(_net_68&_net_78)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))&(_net_68&_net_77)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))&(_net_68&_net_76)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))&(_net_68&_net_75)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))&(_net_68&_net_74)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))&(_net_68&_net_73)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))&(_net_68&_net_72)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))&(_net_68&_net_71)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))&(_net_68&_net_70)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))&(_net_68&_net_69)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))&(_net_35&_net_67)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))&(_net_35&_net_66)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))&(_net_35&_net_65)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))&(_net_35&_net_64)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))&(_net_35&_net_63)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))&(_net_35&_net_62)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))&(_net_35&_net_61)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))&(_net_35&_net_60)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))&(_net_35&_net_59)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))&(_net_35&_net_58)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))&(_net_35&_net_57)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))&(_net_35&_net_56)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))&(_net_35&_net_55)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))&(_net_35&_net_54)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))&(_net_35&_net_53)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))&(_net_35&_net_52)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))&(_net_35&_net_51)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))&(_net_35&_net_50)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))&(_net_35&_net_49)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))&(_net_35&_net_48)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))&(_net_35&_net_47)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))&(_net_35&_net_46)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))&(_net_35&_net_45)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))&(_net_35&_net_44)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))&(_net_35&_net_43)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))&(_net_35&_net_42)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))&(_net_35&_net_41)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))&(_net_35&_net_40)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))&(_net_35&_net_39)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))&(_net_35&_net_38)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))&(_net_35&_net_37)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))&(_net_35&_net_36)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))&(_net_2&_net_34)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))&(_net_2&_net_33)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))&(_net_2&_net_32)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))&(_net_2&_net_31)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))&(_net_2&_net_30)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))&(_net_2&_net_29)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))&(_net_2&_net_28)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))&(_net_2&_net_27)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))&(_net_2&_net_26)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))&(_net_2&_net_25)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))&(_net_2&_net_24)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))&(_net_2&_net_23)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))&(_net_2&_net_22)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))&(_net_2&_net_21)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))&(_net_2&_net_20)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))&(_net_2&_net_19)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))&(_net_2&_net_18)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))&(_net_2&_net_17)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))&(_net_2&_net_16)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))&(_net_2&_net_15)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))&(_net_2&_net_14)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))&(_net_2&_net_13)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))&(_net_2&_net_12)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))&(_net_2&_net_11)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))&(_net_2&_net_10)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))&(_net_2&_net_9)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))&(_net_2&_net_8)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))&(_net_2&_net_7)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))&(_net_2&_net_6)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))|(_net_2&_net_6))&(_net_2&_net_5)))|(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))|(_net_2&_net_6))|(_net_2&_net_5))&(_net_2&_net_4)))|((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))|(_net_2&_net_6))|(_net_2&_net_5))|(_net_2&_net_4))&(_net_2&_net_3))))? 4'bx :(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_net_101&_net_133)|(_net_101&_net_132))|(_net_101&_net_131))|(_net_101&_net_130))|(_net_101&_net_129))|(_net_101&_net_128))|(_net_101&_net_127))|(_net_101&_net_126))|(_net_101&_net_125))|(_net_101&_net_124))|(_net_101&_net_123))|(_net_101&_net_122))|(_net_101&_net_121))|(_net_101&_net_120))|(_net_101&_net_119))|(_net_101&_net_118))|(_net_101&_net_117))|(_net_101&_net_116))|(_net_101&_net_115))|(_net_101&_net_114))|(_net_101&_net_113))|(_net_101&_net_112))|(_net_101&_net_111))|(_net_101&_net_110))|(_net_101&_net_109))|(_net_101&_net_108))|(_net_101&_net_107))|(_net_101&_net_106))|(_net_101&_net_105))|(_net_101&_net_104))|(_net_101&_net_103))|(_net_101&_net_102))|(_net_68&_net_100))|(_net_68&_net_99))|(_net_68&_net_98))|(_net_68&_net_97))|(_net_68&_net_96))|(_net_68&_net_95))|(_net_68&_net_94))|(_net_68&_net_93))|(_net_68&_net_92))|(_net_68&_net_91))|(_net_68&_net_90))|(_net_68&_net_89))|(_net_68&_net_88))|(_net_68&_net_87))|(_net_68&_net_86))|(_net_68&_net_85))|(_net_68&_net_84))|(_net_68&_net_83))|(_net_68&_net_82))|(_net_68&_net_81))|(_net_68&_net_80))|(_net_68&_net_79))|(_net_68&_net_78))|(_net_68&_net_77))|(_net_68&_net_76))|(_net_68&_net_75))|(_net_68&_net_74))|(_net_68&_net_73))|(_net_68&_net_72))|(_net_68&_net_71))|(_net_68&_net_70))|(_net_68&_net_69))|(_net_35&_net_67))|(_net_35&_net_66))|(_net_35&_net_65))|(_net_35&_net_64))|(_net_35&_net_63))|(_net_35&_net_62))|(_net_35&_net_61))|(_net_35&_net_60))|(_net_35&_net_59))|(_net_35&_net_58))|(_net_35&_net_57))|(_net_35&_net_56))|(_net_35&_net_55))|(_net_35&_net_54))|(_net_35&_net_53))|(_net_35&_net_52))|(_net_35&_net_51))|(_net_35&_net_50))|(_net_35&_net_49))|(_net_35&_net_48))|(_net_35&_net_47))|(_net_35&_net_46))|(_net_35&_net_45))|(_net_35&_net_44))|(_net_35&_net_43))|(_net_35&_net_42))|(_net_35&_net_41))|(_net_35&_net_40))|(_net_35&_net_39))|(_net_35&_net_38))|(_net_35&_net_37))|(_net_35&_net_36))|(_net_2&_net_34))|(_net_2&_net_33))|(_net_2&_net_32))|(_net_2&_net_31))|(_net_2&_net_30))|(_net_2&_net_29))|(_net_2&_net_28))|(_net_2&_net_27))|(_net_2&_net_26))|(_net_2&_net_25))|(_net_2&_net_24))|(_net_2&_net_23))|(_net_2&_net_22))|(_net_2&_net_21))|(_net_2&_net_20))|(_net_2&_net_19))|(_net_2&_net_18))|(_net_2&_net_17))|(_net_2&_net_16))|(_net_2&_net_15))|(_net_2&_net_14))|(_net_2&_net_13))|(_net_2&_net_12))|(_net_2&_net_11))|(_net_2&_net_10))|(_net_2&_net_9))|(_net_2&_net_8))|(_net_2&_net_7))|(_net_2&_net_6))|(_net_2&_net_5))|(_net_2&_net_4))|(_net_2&_net_3)))? 
// synthesis translate_on
// synopsys translate_on
(((_net_101&_net_133))?Vin:4'b0)|
    (((_net_101&_net_132))?Vin:4'b0)|
    (((_net_101&_net_131))?Vin:4'b0)|
    (((_net_101&_net_130))?Vin:4'b0)|
    (((_net_101&_net_129))?Vin:4'b0)|
    (((_net_101&_net_128))?Vin:4'b0)|
    (((_net_101&_net_127))?Vin:4'b0)|
    (((_net_101&_net_126))?Vin:4'b0)|
    (((_net_101&_net_125))?Vin:4'b0)|
    (((_net_101&_net_124))?Vin:4'b0)|
    (((_net_101&_net_123))?Vin:4'b0)|
    (((_net_101&_net_122))?Vin:4'b0)|
    (((_net_101&_net_121))?Vin:4'b0)|
    (((_net_101&_net_120))?Vin:4'b0)|
    (((_net_101&_net_119))?Vin:4'b0)|
    (((_net_101&_net_118))?Vin:4'b0)|
    (((_net_101&_net_117))?Vin:4'b0)|
    (((_net_101&_net_116))?Vin:4'b0)|
    (((_net_101&_net_115))?Vin:4'b0)|
    (((_net_101&_net_114))?Vin:4'b0)|
    (((_net_101&_net_113))?Vin:4'b0)|
    (((_net_101&_net_112))?Vin:4'b0)|
    (((_net_101&_net_111))?Vin:4'b0)|
    (((_net_101&_net_110))?Vin:4'b0)|
    (((_net_101&_net_109))?4'b0000:4'b0)|
    (((_net_101&_net_108))?4'b0000:4'b0)|
    (((_net_101&_net_107))?4'b0000:4'b0)|
    (((_net_101&_net_106))?4'b0000:4'b0)|
    (((_net_101&_net_105))?4'b0000:4'b0)|
    (((_net_101&_net_104))?4'b0000:4'b0)|
    (((_net_101&_net_103))?4'b0000:4'b0)|
    (((_net_101&_net_102))?4'b0000:4'b0)|
    (((_net_68&_net_100))?Vin:4'b0)|
    (((_net_68&_net_99))?Vin:4'b0)|
    (((_net_68&_net_98))?Vin:4'b0)|
    (((_net_68&_net_97))?Vin:4'b0)|
    (((_net_68&_net_96))?Vin:4'b0)|
    (((_net_68&_net_95))?Vin:4'b0)|
    (((_net_68&_net_94))?Vin:4'b0)|
    (((_net_68&_net_93))?Vin:4'b0)|
    (((_net_68&_net_92))?Vin:4'b0)|
    (((_net_68&_net_91))?Vin:4'b0)|
    (((_net_68&_net_90))?Vin:4'b0)|
    (((_net_68&_net_89))?Vin:4'b0)|
    (((_net_68&_net_88))?Vin:4'b0)|
    (((_net_68&_net_87))?Vin:4'b0)|
    (((_net_68&_net_86))?Vin:4'b0)|
    (((_net_68&_net_85))?Vin:4'b0)|
    (((_net_68&_net_84))?4'b0000:4'b0)|
    (((_net_68&_net_83))?4'b0000:4'b0)|
    (((_net_68&_net_82))?4'b0000:4'b0)|
    (((_net_68&_net_81))?4'b0000:4'b0)|
    (((_net_68&_net_80))?4'b0000:4'b0)|
    (((_net_68&_net_79))?4'b0000:4'b0)|
    (((_net_68&_net_78))?4'b0000:4'b0)|
    (((_net_68&_net_77))?4'b0000:4'b0)|
    (((_net_68&_net_76))?4'b0000:4'b0)|
    (((_net_68&_net_75))?4'b0000:4'b0)|
    (((_net_68&_net_74))?4'b0000:4'b0)|
    (((_net_68&_net_73))?4'b0000:4'b0)|
    (((_net_68&_net_72))?4'b0000:4'b0)|
    (((_net_68&_net_71))?4'b0000:4'b0)|
    (((_net_68&_net_70))?4'b0000:4'b0)|
    (((_net_68&_net_69))?4'b0000:4'b0)|
    (((_net_35&_net_67))?Vin:4'b0)|
    (((_net_35&_net_66))?Vin:4'b0)|
    (((_net_35&_net_65))?Vin:4'b0)|
    (((_net_35&_net_64))?Vin:4'b0)|
    (((_net_35&_net_63))?Vin:4'b0)|
    (((_net_35&_net_62))?Vin:4'b0)|
    (((_net_35&_net_61))?Vin:4'b0)|
    (((_net_35&_net_60))?Vin:4'b0)|
    (((_net_35&_net_59))?4'b0000:4'b0)|
    (((_net_35&_net_58))?4'b0000:4'b0)|
    (((_net_35&_net_57))?4'b0000:4'b0)|
    (((_net_35&_net_56))?4'b0000:4'b0)|
    (((_net_35&_net_55))?4'b0000:4'b0)|
    (((_net_35&_net_54))?4'b0000:4'b0)|
    (((_net_35&_net_53))?4'b0000:4'b0)|
    (((_net_35&_net_52))?4'b0000:4'b0)|
    (((_net_35&_net_51))?4'b0000:4'b0)|
    (((_net_35&_net_50))?4'b0000:4'b0)|
    (((_net_35&_net_49))?4'b0000:4'b0)|
    (((_net_35&_net_48))?4'b0000:4'b0)|
    (((_net_35&_net_47))?4'b0000:4'b0)|
    (((_net_35&_net_46))?4'b0000:4'b0)|
    (((_net_35&_net_45))?4'b0000:4'b0)|
    (((_net_35&_net_44))?4'b0000:4'b0)|
    (((_net_35&_net_43))?4'b0000:4'b0)|
    (((_net_35&_net_42))?4'b0000:4'b0)|
    (((_net_35&_net_41))?4'b0000:4'b0)|
    (((_net_35&_net_40))?4'b0000:4'b0)|
    (((_net_35&_net_39))?4'b0000:4'b0)|
    (((_net_35&_net_38))?4'b0000:4'b0)|
    (((_net_35&_net_37))?4'b0000:4'b0)|
    (((_net_35&_net_36))?4'b0000:4'b0)|
    (((_net_2&_net_34))?Vin:4'b0)|
    (((_net_2&_net_33))?Vin:4'b0)|
    (((_net_2&_net_32))?Vin:4'b0)|
    (((_net_2&_net_31))?Vin:4'b0)|
    (((_net_2&_net_30))?4'b0000:4'b0)|
    (((_net_2&_net_29))?4'b0000:4'b0)|
    (((_net_2&_net_28))?4'b0000:4'b0)|
    (((_net_2&_net_27))?4'b0000:4'b0)|
    (((_net_2&_net_26))?4'b0000:4'b0)|
    (((_net_2&_net_25))?4'b0000:4'b0)|
    (((_net_2&_net_24))?4'b0000:4'b0)|
    (((_net_2&_net_23))?4'b0000:4'b0)|
    (((_net_2&_net_22))?4'b0000:4'b0)|
    (((_net_2&_net_21))?4'b0000:4'b0)|
    (((_net_2&_net_20))?4'b0000:4'b0)|
    (((_net_2&_net_19))?4'b0000:4'b0)|
    (((_net_2&_net_18))?4'b0000:4'b0)|
    (((_net_2&_net_17))?4'b0000:4'b0)|
    (((_net_2&_net_16))?4'b0000:4'b0)|
    (((_net_2&_net_15))?4'b0000:4'b0)|
    (((_net_2&_net_14))?4'b0000:4'b0)|
    (((_net_2&_net_13))?4'b0000:4'b0)|
    (((_net_2&_net_12))?4'b0000:4'b0)|
    (((_net_2&_net_11))?4'b0000:4'b0)|
    (((_net_2&_net_10))?4'b0000:4'b0)|
    (((_net_2&_net_9))?4'b0000:4'b0)|
    (((_net_2&_net_8))?4'b0000:4'b0)|
    (((_net_2&_net_7))?4'b0000:4'b0)|
    (((_net_2&_net_6))?4'b0000:4'b0)|
    (((_net_2&_net_5))?4'b0000:4'b0)|
    (((_net_2&_net_4))?4'b0000:4'b0)|
    (((_net_2&_net_3))?4'b0000:4'b0)
// synthesis translate_off
// synopsys translate_off
:4'bx
// synthesis translate_on
// synopsys translate_on
;
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     cnt <= 6'b000000;
else 
// synthesis translate_off
// synopsys translate_off
if ((((exec&_net_1)&(exec&_net_0))|(((exec&_net_1)|(exec&_net_0))&setduty)))   cnt <= 6'bx; 
  else 
// synthesis translate_on
// synopsys translate_on
if ((exec&_net_1))
      cnt <= 6'b000000;
else if ((exec&_net_0))
      cnt <= (cnt+6'b000001);
else if (setduty)
      cnt <= 6'b000000;
end

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock)
  begin
if (((((exec&_net_1)|(exec&_net_0))|setduty)==1'b1) ||
 ((((exec&_net_1)|(exec&_net_0))|setduty)==1'b0) ) begin
 if ((((exec&_net_1)&(exec&_net_0))|(((exec&_net_1)|(exec&_net_0))&setduty)))
 begin $display("Warning: assign collision(duty2:cnt) at %d",$time);

  end
 end
 else 
 $display("Warning: register set hazard(duty2:cnt) at %d",$time);

  end

// synthesis translate_on
// synopsys translate_on
always @(posedge m_clock)
  begin
if (setduty)
      d <= dnum;
end
endmodule
/*
 Produced by NSL Core(version=20140126), IP ARCH, Inc. Sun Aug 14 20:41:11 2016
 Licensed to :EVALUATION USER
*/
